library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity rom_char_l is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of rom_char_l is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"04",X"0C",X"02",X"02",X"FE",X"FE",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"26",X"AF",X"AF",X"AF",X"2E",X"FC",X"00",X"0F",X"FE",X"16",X"0E",X"16",X"FE",X"0F",X"00",
		X"68",X"FA",X"9B",X"0B",X"9B",X"FA",X"68",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",
		X"10",X"10",X"10",X"FF",X"FF",X"10",X"10",X"10",X"00",X"E7",X"A5",X"E5",X"E5",X"A5",X"E7",X"00",
		X"3F",X"63",X"41",X"00",X"00",X"41",X"63",X"3F",X"00",X"30",X"20",X"20",X"20",X"20",X"20",X"00",
		X"00",X"70",X"50",X"40",X"70",X"10",X"70",X"00",X"00",X"70",X"40",X"70",X"40",X"40",X"70",X"00",
		X"00",X"10",X"10",X"50",X"50",X"70",X"40",X"00",X"00",X"70",X"10",X"70",X"40",X"40",X"70",X"00",
		X"00",X"70",X"10",X"70",X"50",X"50",X"70",X"00",X"00",X"70",X"40",X"40",X"40",X"40",X"40",X"00",
		X"00",X"70",X"50",X"70",X"50",X"50",X"70",X"00",X"00",X"70",X"50",X"70",X"40",X"40",X"40",X"00",
		X"00",X"00",X"00",X"80",X"C0",X"E0",X"F0",X"F8",X"00",X"04",X"0F",X"FF",X"FB",X"E5",X"9E",X"6E",
		X"00",X"0F",X"B7",X"57",X"DB",X"CB",X"9C",X"9C",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"13",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"D8",
		X"00",X"00",X"00",X"00",X"00",X"80",X"E0",X"F8",X"00",X"00",X"00",X"00",X"04",X"0D",X"13",X"9F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"BC",X"BF",X"BC",X"BC",X"BC",
		X"00",X"00",X"00",X"01",X"07",X"01",X"01",X"81",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"0D",
		X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"3C",X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"1C",
		X"00",X"18",X"6C",X"EE",X"6C",X"6C",X"6C",X"6C",X"00",X"00",X"00",X"10",X"DC",X"B0",X"30",X"D8",
		X"FC",X"F0",X"C6",X"88",X"60",X"80",X"00",X"00",X"01",X"03",X"0F",X"3F",X"FC",X"F1",X"E6",X"9C",
		X"9C",X"9C",X"8C",X"88",X"80",X"83",X"87",X"8F",X"DD",X"9D",X"89",X"8B",X"97",X"95",X"B5",X"A9",
		X"1D",X"1D",X"0D",X"0D",X"0D",X"0D",X"F1",X"8D",X"DE",X"B2",X"B6",X"B5",X"AF",X"A7",X"66",X"07",
		X"F0",X"70",X"60",X"61",X"61",X"61",X"61",X"61",X"AC",X"AF",X"AF",X"A3",X"A3",X"A3",X"A3",X"B3",
		X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"0D",X"BC",X"BC",X"BC",X"BC",X"BC",X"BC",X"BC",X"7C",
		X"E1",X"11",X"71",X"71",X"71",X"71",X"6E",X"71",X"0D",X"8B",X"8B",X"9B",X"9A",X"9A",X"96",X"94",
		X"DF",X"EF",X"F7",X"7B",X"3B",X"1B",X"1B",X"1B",X"DB",X"EB",X"E0",X"60",X"60",X"60",X"20",X"20",
		X"6C",X"6C",X"6C",X"AC",X"5C",X"3C",X"DC",X"EC",X"EC",X"F4",X"7C",X"3F",X"1C",X"1D",X"15",X"11",
		X"30",X"F8",X"FC",X"FC",X"0E",X"76",X"F6",X"3C",X"20",X"01",X"03",X"07",X"1F",X"FE",X"F8",X"F2",
		X"AF",X"AF",X"AF",X"AF",X"AF",X"B7",X"D3",X"19",X"AD",X"CD",X"FD",X"DD",X"AD",X"8D",X"8D",X"0C",
		X"1D",X"8D",X"CD",X"CD",X"AD",X"ED",X"E9",X"80",X"43",X"C6",X"FC",X"D3",X"9D",X"B1",X"80",X"00",
		X"63",X"62",X"62",X"66",X"66",X"65",X"75",X"00",X"D3",X"61",X"61",X"B3",X"BB",X"C3",X"C3",X"C2",
		X"26",X"6B",X"7D",X"5D",X"0E",X"0E",X"05",X"03",X"BC",X"BC",X"BC",X"BC",X"BC",X"BC",X"9C",X"EE",
		X"39",X"4B",X"DB",X"39",X"B5",X"3D",X"1D",X"10",X"B4",X"AC",X"2F",X"6D",X"69",X"5B",X"5C",X"80",
		X"17",X"17",X"37",X"2F",X"1E",X"FE",X"F8",X"00",X"00",X"00",X"00",X"00",X"88",X"A7",X"79",X"3E",
		X"EC",X"6C",X"6C",X"6E",X"9F",X"3F",X"CC",X"F1",X"28",X"28",X"2C",X"5E",X"B9",X"DA",X"EB",X"F1",
		X"3C",X"18",X"10",X"10",X"20",X"00",X"60",X"C0",X"F4",X"40",X"40",X"80",X"80",X"00",X"00",X"00",
		X"BC",X"9E",X"0F",X"07",X"03",X"01",X"00",X"00",X"0F",X"8F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C1",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"C3",X"87",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"9F",X"FF",X"FF",X"FC",X"70",X"00",X"B8",X"F7",X"7B",X"3D",X"1E",X"0E",X"07",X"07",X"03",
		X"19",X"3C",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"E1",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"07",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"20",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"FF",X"00",X"00",X"00",X"00",X"F0",X"FF",X"FF",X"FF",
		X"00",X"00",X"F8",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"0F",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"FC",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FC",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"FC",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"3F",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"3F",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"3F",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"FF",X"00",X"00",X"00",X"00",X"00",X"F0",X"FF",X"FF",
		X"00",X"00",X"80",X"F0",X"FF",X"FF",X"FF",X"FF",X"F8",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"C0",X"F8",X"FF",X"FF",
		X"00",X"00",X"80",X"FC",X"FF",X"FF",X"FF",X"FF",X"00",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F8",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"1F",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"03",X"1F",X"FF",X"FF",X"1F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"00",X"01",X"0F",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"FF",X"00",X"00",X"00",X"00",X"C0",X"F8",X"FF",X"FF",
		X"80",X"E0",X"F8",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"80",X"E0",X"F8",X"FE",X"80",X"E0",X"F8",X"FE",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"80",X"E0",X"F8",X"FF",
		X"00",X"00",X"F0",X"FE",X"FF",X"FF",X"FF",X"FF",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"07",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"0F",X"7F",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"07",X"1F",X"7F",
		X"01",X"07",X"1F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"01",X"07",X"1F",X"7F",X"01",X"07",X"1F",X"7F",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"03",X"1F",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"FF",X"00",X"00",X"C0",X"F0",X"FC",X"FF",X"FF",X"FF",
		X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"80",X"C0",X"F0",X"F8",
		X"F0",X"F8",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",
		X"00",X"C0",X"E0",X"F0",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"F8",X"FE",X"00",X"80",X"F0",X"FC",X"FF",X"FF",X"FF",X"FF",
		X"F8",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"01",X"0F",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"07",X"1F",X"7F",X"00",X"03",X"07",X"0F",X"3F",X"FF",X"FF",X"FF",
		X"0F",X"1F",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",
		X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"03",X"0F",X"1F",
		X"00",X"00",X"03",X"0F",X"3F",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"00",X"33",X"33",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"FF",X"00",X"C0",X"E0",X"F0",X"F8",X"FE",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"80",X"E0",X"F0",X"F8",X"FC",X"FE",
		X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"80",X"C0",X"E0",X"E0",X"F0",X"F8",X"FC",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"80",X"80",X"C0",X"E0",X"F0",X"F8",X"FC",X"FE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"80",X"E0",X"F0",X"F8",X"FC",X"FE",X"FF",
		X"3E",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"07",X"0F",X"3F",X"FF",X"FF",
		X"03",X"0F",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"E0",X"F0",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"1E",X"7F",X"FF",
		X"03",X"0F",X"1F",X"3F",X"7F",X"FF",X"FF",X"FF",X"07",X"0F",X"1F",X"3F",X"7F",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"0F",X"1F",X"3F",X"7F",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"0F",X"1F",X"3F",X"7F",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"F8",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"1F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"F8",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"1F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"80",X"C0",X"F8",X"FF",X"E0",X"F8",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"F0",X"F8",X"FC",X"FE",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"F8",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"80",X"C0",X"C0",X"E0",X"F0",X"F8",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"C0",X"E0",X"F0",X"F8",X"F8",X"FC",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"F0",X"F0",X"FC",X"FC",X"FE",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"80",X"80",X"C0",X"E0",X"F0",
		X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"80",X"C0",X"C0",X"E0",X"F0",X"F8",X"F8",X"FC",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"F8",X"FC",X"FE",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"1F",X"3F",X"7F",X"FF",
		X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"01",X"03",X"03",X"07",X"0F",X"0F",X"1F",X"3F",
		X"0F",X"1F",X"3F",X"3F",X"7F",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"0F",
		X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"03",X"03",X"07",X"0F",X"1F",X"1F",X"3F",X"7F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"1F",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"01",X"03",X"03",X"07",X"0F",X"1F",X"07",X"0F",X"1F",X"3F",X"7F",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"07",X"0F",X"1F",X"3F",X"7F",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"00",X"00",X"00",X"00",X"00",X"01",X"1F",X"FF",
		X"FF",X"F8",X"E0",X"C0",X"80",X"80",X"00",X"00",X"C0",X"C0",X"80",X"80",X"80",X"80",X"00",X"00",
		X"F0",X"F0",X"E0",X"E0",X"E0",X"E0",X"C0",X"C0",X"F8",X"F8",X"F8",X"F8",X"F0",X"F0",X"F0",X"F0",
		X"FE",X"FE",X"FE",X"FE",X"FC",X"FC",X"FC",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"E0",X"E0",X"E0",X"C0",X"C0",X"C0",
		X"FC",X"FC",X"FC",X"F8",X"F8",X"F8",X"F8",X"F0",X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",X"FE",X"FC",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"F8",X"E0",X"C0",
		X"FF",X"FF",X"FF",X"7F",X"3F",X"1F",X"07",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"07",X"07",X"03",X"03",X"03",X"01",X"01",X"1F",X"1F",X"1F",X"0F",X"0F",X"0F",X"0F",X"07",
		X"7F",X"7F",X"7F",X"3F",X"3F",X"3F",X"3F",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"03",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"0F",X"07",X"07",X"07",X"07",X"03",X"03",X"03",
		X"1F",X"1F",X"1F",X"1F",X"0F",X"0F",X"0F",X"0F",X"7F",X"7F",X"7F",X"7F",X"3F",X"3F",X"3F",X"3F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"07",X"03",X"01",X"01",X"00",X"00",
		X"FF",X"FC",X"F8",X"F0",X"E0",X"C0",X"C0",X"80",X"F0",X"E0",X"C0",X"C0",X"80",X"80",X"00",X"00",
		X"FF",X"FF",X"FE",X"FE",X"FC",X"FC",X"F8",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FE",X"FC",X"F8",X"F8",X"F8",X"F0",X"E0",X"C0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",
		X"1F",X"1F",X"0F",X"0F",X"07",X"03",X"03",X"01",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"3F",
		X"FF",X"F7",X"E1",X"C1",X"C0",X"80",X"00",X"00",X"7C",X"38",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"0F",X"07",X"07",X"03",X"03",X"01",X"01",X"00",
		X"FF",X"FF",X"FF",X"7F",X"3F",X"3F",X"1F",X"1F",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"1F",X"0F",X"07",X"07",X"03",X"03",X"01",X"FF",X"F8",X"F0",X"E0",X"C0",X"80",X"00",X"00",
		X"FC",X"F8",X"F0",X"E0",X"C0",X"80",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",
		X"FC",X"F8",X"70",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",
		X"FF",X"F1",X"C0",X"80",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"78",
		X"3F",X"1F",X"0F",X"07",X"03",X"01",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",
		X"1F",X"0F",X"07",X"03",X"01",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",X"3F",
		X"FF",X"1F",X"07",X"01",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"00",
		X"E0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"80",X"F0",X"F0",X"F0",X"E0",X"E0",X"E0",X"E0",X"E0",
		X"FF",X"FE",X"FC",X"FC",X"F8",X"F8",X"F8",X"F0",X"FC",X"FC",X"F8",X"F8",X"F0",X"F0",X"E0",X"C0",
		X"FF",X"FF",X"FE",X"FE",X"FE",X"FE",X"FE",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3F",X"1F",X"1F",X"1F",X"0F",X"0F",X"07",X"03",X"FF",X"FF",X"7F",X"7F",X"7D",X"7D",X"3F",X"3F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",
		X"07",X"03",X"03",X"03",X"03",X"03",X"03",X"01",X"0F",X"0F",X"0F",X"07",X"07",X"07",X"07",X"07",
		X"FF",X"7F",X"3F",X"3F",X"1F",X"1F",X"1F",X"0F",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",
		X"FF",X"FC",X"F0",X"F0",X"E0",X"C0",X"C0",X"C0",X"FC",X"FC",X"F8",X"F8",X"F0",X"F0",X"E0",X"C0",
		X"FF",X"FE",X"FE",X"FE",X"FE",X"FE",X"FC",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3F",X"3F",X"1F",X"1F",X"0F",X"0F",X"07",X"03",X"FF",X"7F",X"7F",X"7F",X"7F",X"7F",X"3F",X"3F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",
		X"FF",X"3F",X"0F",X"0F",X"07",X"03",X"03",X"03",X"00",X"00",X"00",X"00",X"C0",X"F0",X"FC",X"FF",
		X"C0",X"F0",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"C0",X"F0",X"FC",X"FF",X"C0",X"F0",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"C0",X"F0",X"FC",X"FF",
		X"C0",X"F0",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"C0",X"F0",X"FC",X"FF",X"C0",X"F0",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"E7",X"F7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"FF",X"FF",X"FF",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"07",X"07",X"07",X"03",X"03",X"03",X"01",X"00",X"FF",X"FF",X"7F",X"3F",X"1F",X"1F",X"0F",X"0F",
		X"E3",X"E3",X"E3",X"E3",X"E3",X"E3",X"F3",X"FB",X"FF",X"FF",X"FF",X"FF",X"E3",X"E3",X"E3",X"E3",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F9",X"FD",X"FF",X"FF",X"3F",X"0F",X"07",X"03",X"FF",X"FF",X"FF",X"FF",X"F1",X"F1",X"F1",X"F1",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"3F",X"07",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"38",X"38",X"FC",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FC",X"E0",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"1C",X"1C",X"3F",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"9F",X"BF",X"FF",X"FF",X"FC",X"F0",X"E0",X"C0",X"FF",X"FF",X"FF",X"FF",X"8F",X"8F",X"8F",X"8F",
		X"E0",X"E0",X"E0",X"C0",X"C0",X"C0",X"80",X"80",X"FF",X"FF",X"FE",X"FC",X"F8",X"F8",X"F0",X"F0",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"CF",X"DF",X"FF",X"FF",X"FF",X"FF",X"C7",X"C7",X"C7",X"C7",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E3",X"E3",X"E3",X"E3",X"E3",X"E3",X"E7",X"EF",
		X"E3",X"E3",X"E3",X"E3",X"E3",X"E3",X"E3",X"E3",X"FF",X"FF",X"FF",X"FF",X"E3",X"E3",X"E3",X"E3",
		X"03",X"0F",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"03",X"0F",X"3F",X"FF",X"03",X"0F",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"03",X"0F",X"3F",X"FF",
		X"03",X"0F",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"03",X"0F",X"3F",X"FF",X"03",X"0F",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"03",X"0F",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
